module binary_bcd_2(bin_in, digit_1, digit_2);
  
  input [6:0] bin_in;
  output [3:0] digit_1;
  output [3:0] digit_2;
  
  // Binary-to-BCD logic goes here
  
endmodule